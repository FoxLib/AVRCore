
// Заполнение данными регистров
// ---------------------------------------------------------------------

initial begin

    // Выводы
    we = 0; o_data = 0; pc = 0; address = 0;

    // Регистры 0-15
    r[0] = 8'h00; r[4] = 8'h00; r[8]  = 8'h00; r[12] = 8'h01;
    r[1] = 8'h00; r[5] = 8'h00; r[9]  = 8'h00; r[13] = 8'h00;
    r[2] = 8'h00; r[6] = 8'h00; r[10] = 8'h00; r[14] = 8'h00;
    r[3] = 8'h00; r[7] = 8'h00; r[11] = 8'h00; r[15] = 8'h00;

    // Регистры 16-31
    r[16] = 8'h00; r[20] = 8'h00; r[24] = 8'h00; r[28] = 8'h00;
    r[17] = 8'h00; r[21] = 8'h00; r[25] = 8'h00; r[29] = 8'h00;
    r[18] = 8'h00; r[22] = 8'h00; r[26] = 8'h00; r[30] = 8'h05;
    r[19] = 8'h00; r[23] = 8'h00; r[27] = 8'h00; r[31] = 8'hFA;

end


// Проксирование памяти
// ---------------------------------------------------------------------

always @* begin

    casex (address)

        // Регистры
        16'b0000_0000_000x_xxxx: din = r[ address[4:0] ];

        // Процессор
        16'h005B: din = rampz;
        16'h005D: din = sp[ 7:0];
        16'h005E: din = sp[15:8];
        16'h005F: din = sreg;

        // Память
        default:  din = i_data;

    endcase

end

// Текущее состояние процессора
// ---------------------------------------------------------------------
reg [ 7:0]  din;
reg [ 7:0]  rampz   = 0;
reg [ 3:0]  st      = 0;            // Машина состояний
reg [ 3:0]  stnext  = 0;            // Следующий код состояния
reg [ 7:0]  latch   = 0;            // Защелка опкода
reg [ 7:0]  r[32];                  // Регистры
reg [15:0]  sp;                     // Стек
reg [ 7:0]  sreg;                   // Флаги

// Управление
// ---------------------------------------------------------------------
reg         pcload;                 // =1 Загрузка из pcnext
reg [15:0]  pcnext;
reg         reg_w;                  // =1 Запись АЛУ в регистр reg_id
reg         sreg_w;                 // =1 Запись из АЛУ в регистр флагов
reg [ 4:0]  reg_id;                 // Номер регистра
reg         wren;                   // Запись в память
reg [ 7:0]  wdata;

// Провода
// ---------------------------------------------------------------------
wire [15:0] opcode = st ? latch : ir;
wire [15:0] X   = {r[27], r[26]};
wire [15:0] Y   = {r[29], r[28]};
wire [15:0] Z   = {r[31], r[30]};
wire [15:0] Xm  = X - 1;
wire [15:0] Xp  = X + 1;
wire [15:0] Ym  = Y - 1;
wire [15:0] Yp  = Y + 1;
wire [15:0] Zm  = Z - 1;
wire [15:0] Zp  = Z + 1;
wire [ 5:0] q   = {opcode[13], opcode[11:10], opcode[2:0]};
wire [ 4:0] rd  =  opcode[8:4];
wire [ 4:0] rr  = {opcode[9], opcode[3:0]};
wire [ 4:0] rdi = {1'b1, opcode[7:4]};
wire [ 4:0] rri = {1'b1, opcode[3:0]};
wire [ 7:0] K   = {opcode[11:8], opcode[3:0]};
