`timescale 10ns / 1ns

module avr;

// ---------------------------------------------------------------------
// Симулятор Verilog Icarus
// ---------------------------------------------------------------------

reg clock  = 0;
reg clk50  = 0;
reg clklo  = 0;
reg locked = 0;

always #0.5 clock = ~clock;
always #1.0 clk50 = ~clk50;
always #1.5 clklo = ~clklo;

initial begin clock = 0; clk50 = 1; clklo = 0; #3.0 locked = 1; #2000 $finish; end
initial begin $dumpfile("tb.vcd"); $dumpvars(0, avr); end

// ---------------------------------------------------------------------
// Интерфейс для работы с памятью (чтение и запись)
// ---------------------------------------------------------------------

reg [15:0] flash[ 65536]; // 128k
reg [ 7:0] sram [131072]; // 128k

initial $readmemh("mem_core.hex", flash, 16'h0000);
initial $readmemh("mem_sram.hex", sram,  16'h0000);

// ---------------------------------------------------------------------
// Основной интерфейс ядра
// ---------------------------------------------------------------------

wire [15:0] pc;         // Программный счетчик
reg  [15:0] ir;         // Регистр инструкции (текущий опкод)
wire [15:0] address;    // Адрес в память SRAM
reg  [ 7:0] data_i;     // Прочтенные данные из SRAM
wire [ 7:0] data_o;     // Данные для записи в SRAM
wire [ 7:0] wren;       // Разрешение на запись в память

// Контроллер внутрисхемной памяти
always @(posedge clock) begin

    ir     <= flash[     pc];
    data_i <= sram [address];

    if (wren) sram[address] <= data_o;

end

// ---------------------------------------------------------------------
// Центральный процессорный блок
// ---------------------------------------------------------------------

/*
cpu UnitAVRCPU
(
    // Тактовый генератор
    .clock      (clklo & locked),

    // Программная память
    .pc         (pc),          // Программный счетчик
    .ir         (ir),          // Инструкция из памяти

    // Оперативная память
    .address    (mem_ad),       // Указатель на память RAM (sram)
    .din        (mem),          // memory[ address ]
    .wb         (mem_wb),       // Запись в память по address
    .w          (mem_w),        // Разрешение записи в память
);
*/

endmodule
